

module mul_l3(W1234,W5678,W9101112,W13141516,W17181920,W21222324,OUT12345678,OUT910111213141516,OUT1718192021222324);
		
        input  [5:0]  W1234;
		input  [9:0]  W5678;
		input  [13:0] W9101112;
		input  [17:0] W13141516;
		input  [21:0] W17181920;
		input  [24:0] W21222324;
		output [10:0] OUT12345678;
		output [18:0] OUT910111213141516;
		output [24:0] OUT1718192021222324;
	
	
	// LINE 1234, 5678
	wire CARRY12345678_0, CARRY12345678_1;
	cla  l3_00(.A(W1234[3:0]), .B(W5678[3:0]), .CIN(1'b0), .COUT(CARRY12345678_0), .S(OUT12345678[3:0]));
	cla  l3_01(.A({2'b0,W1234[5:4]}), .B(W5678[7:4]), .CIN(CARRY12345678_0), .COUT(CARRY12345678_1), .S(OUT12345678[7:4]));
	tcla l3_02(.A(W5678[9:8]), .CIN(CARRY12345678_1), .COUT(OUT12345678[10]), .S(OUT12345678[9:8]));
	
	// line 9101112, 13141516
	wire CARRY910111213141516_0, CARRY910111213141516_1, CARRY910111213141516_2, CARRY910111213141516_3;
	cla  l3_10(.A(W9101112[3:0]), .B(W13141516[3:0]), .CIN(1'b0), .COUT(CARRY910111213141516_0), .S(OUT910111213141516[3:0]));
	cla  l3_11(.A(W9101112[7:4]), .B(W13141516[7:4]), .CIN(CARRY910111213141516_0), .COUT(CARRY910111213141516_1), .S(OUT910111213141516[7:4]));
	cla  l3_12(.A(W9101112[11:8]), .B(W13141516[11:8]), .CIN(CARRY910111213141516_1), .COUT(CARRY910111213141516_2), .S(OUT910111213141516[11:8]));
	cla  l3_13(.A({2'b0,W9101112[13:12]}), .B(W13141516[15:12]), .CIN(CARRY910111213141516_2), .COUT(CARRY910111213141516_3), .S(OUT910111213141516[15:12]));
	tcla l3_14(.A(W13141516[17:16]), .CIN(CARRY910111213141516_3), .COUT(OUT910111213141516[18]), .S(OUT910111213141516[17:16]));
	
	// line 17181920, 21222324
	wire CARRY1718192021222324_0, CARRY1718192021222324_1, CARRY1718192021222324_2, CARRY1718192021222324_3, CARRY1718192021222324_4, CARRY1718192021222324_5;
	cla l3_20(.A(W17181920[3:0]), .B(W21222324[3:0]), .CIN(1'b0), .COUT(CARRY1718192021222324_0), .S(OUT1718192021222324[3:0]));
	cla l3_21(.A(W17181920[7:4]), .B(W21222324[7:4]), .CIN(CARRY1718192021222324_0), .COUT(CARRY1718192021222324_1), .S(OUT1718192021222324[7:4]));
	cla l3_22(.A(W17181920[11:8]), .B(W21222324[11:8]), .CIN(CARRY1718192021222324_1), .COUT(CARRY1718192021222324_2), .S(OUT1718192021222324[11:8]));
	cla l3_23(.A(W17181920[15:12]), .B(W21222324[15:12]), .CIN(CARRY1718192021222324_2), .COUT(CARRY1718192021222324_3), .S(OUT1718192021222324[15:12]));
	cla l3_24(.A(W17181920[19:16]), .B(W21222324[19:16]), .CIN(CARRY1718192021222324_3), .COUT(CARRY1718192021222324_4), .S(OUT1718192021222324[19:16]));
	cla l3_25(.A({2'b0,W17181920[21:20]}), .B(W21222324[23:20]), .CIN(CARRY1718192021222324_4), .COUT(CARRY1718192021222324_5), .S(OUT1718192021222324[23:20]));
	ha  l3_26(.A(W21222324[24]), .B(CARRY1718192021222324_5), .COUT(), .SUM(OUT1718192021222324[24]));
	
endmodule 

