



module mul_l4(W12345678,W910111213141516,W1718192021222324,OUT12345678910111213141516,OUT1718192021222324);
		input  [10:0] W12345678;
		input  [18:0] W910111213141516;
		input  [24:0] W1718192021222324;
		output [19:0] OUT12345678910111213141516;
		output [24:0] OUT1718192021222324;
	
	
	// line 17181920, 21222324
	wire CARRY12345678910111213141516_0, CARRY12345678910111213141516_1, CARRY12345678910111213141516_2, CARRY12345678910111213141516_3;
	cla  l4_00(.A(W12345678[3:0]), .B(W910111213141516[3:0]), .CIN(1'b0), .COUT(CARRY12345678910111213141516_0), .S(OUT12345678910111213141516[3:0]));
	cla  l4_01(.A(W12345678[7:4]), .B(W910111213141516[7:4]), .CIN(CARRY12345678910111213141516_0), .COUT(CARRY12345678910111213141516_1), .S(OUT12345678910111213141516[7:4]));
	cla  l4_02(.A({1'b0,W12345678[10:8]}), .B(W910111213141516[11:8]), .CIN(CARRY12345678910111213141516_1), .COUT(CARRY12345678910111213141516_2), .S(OUT12345678910111213141516[11:8]));
	ocla l4_03(.A(W910111213141516[15:12]), .CIN(CARRY12345678910111213141516_2), .COUT(CARRY12345678910111213141516_3), .S(OUT12345678910111213141516[15:12]));
	ocla l4_04(.A({1'b0,W910111213141516[18:16]}), .CIN(CARRY12345678910111213141516_3), .COUT(), .S(OUT12345678910111213141516[19:16]));
	
	assign OUT1718192021222324 = W1718192021222324;
	
endmodule 
