



module mul_l2(W12,W34,W56,W78,W910,W1112,W1314,W1516,W1718,W1920,W2122,W2324,OUT1234,OUT5678,OUT9101112,OUT13141516,OUT17181920,OUT21222324);
		
    input  [2:0]  W12;
	input  [4:0]  W34;
	input  [6:0]  W56;
	input  [8:0]  W78;
	input  [10:0] W910;
	input  [12:0] W1112;
	input  [14:0] W1314;
	input  [16:0] W1516;
	input  [18:0] W1718;
	input  [20:0] W1920;
	input  [22:0] W2122;
	input  [24:0] W2324;
	output [5:0]  OUT1234;
	output [9:0]  OUT5678;
	output [13:0] OUT9101112;
	output [17:0] OUT13141516;
	output [21:0] OUT17181920;
	output [24:0] OUT21222324 ;

		
	// line 12, 34
	wire CARRY1234_0;
	cla l2_00(.A({1'b0,W12}), .B(W34[3:0]), .CIN(1'b0), .COUT(CARRY1234_0), .S(OUT1234[3:0]));
	ha  l2_01(.A(W34[4]), .B(CARRY1234_0), .COUT(OUT1234[5]), .SUM(OUT1234[4]));
	
	// line 56, 78
	wire CARRY5678_0, CARRY5678_1;
	cla l2_10(.A(W56[3:0]), .B(W78[3:0]), .CIN(1'b0), .COUT(CARRY5678_0), .S(OUT5678[3:0]));
	cla l2_11(.A({1'b0,W56[6:4]}), .B(W78[7:4]), .CIN(CARRY5678_0), .COUT(CARRY5678_1), .S(OUT5678[7:4]));
	ha  l2_12(.A(W78[8]), .B(CARRY5678_1), .COUT(OUT5678[9]), .SUM(OUT5678[8]));
	
	// line 910, 1112
	wire CARRY9101112_0, CARRY9101112_1, CARRY9101112_2;
	cla l2_20(.A(W910[3:0]), .B(W1112[3:0]), .CIN(1'b0), .COUT(CARRY9101112_0), .S(OUT9101112[3:0]));
	cla l2_21(.A(W910[7:4]), .B(W1112[7:4]), .CIN(CARRY9101112_0), .COUT(CARRY9101112_1), .S(OUT9101112[7:4]));
	cla l2_22(.A({1'b0,W910[10:8]}), .B(W1112[11:8]), .CIN(CARRY9101112_1), .COUT(CARRY9101112_2), .S(OUT9101112[11:8]));
	ha  l2_23(.A(W1112[12]), .B(CARRY9101112_2), .COUT(OUT9101112[13]), .SUM(OUT9101112[12]));
	
	// LINE 1314, 1516
	wire CARRY13141516_0, CARRY13141516_1, CARRY13141516_2, CARRY13141516_3;
	cla l2_30(.A(W1314[3:0]), .B(W1516[3:0]), .CIN(1'b0), .COUT(CARRY13141516_0), .S(OUT13141516[3:0]));
	cla l2_31(.A(W1314[7:4]), .B(W1516[7:4]), .CIN(CARRY13141516_0), .COUT(CARRY13141516_1), .S(OUT13141516[7:4]));
	cla l2_32(.A(W1314[11:8]), .B(W1516[11:8]), .CIN(CARRY13141516_1), .COUT(CARRY13141516_2), .S(OUT13141516[11:8]));
	cla l2_33(.A({1'b0,W1314[14:12]}), .B(W1516[15:12]), .CIN(CARRY13141516_2), .COUT(CARRY13141516_3), .S(OUT13141516[15:12]));
	ha  l2_34(.A(W1516[16]), .B(CARRY13141516_3), .COUT(OUT13141516[17]), .SUM(OUT13141516[16]));
	
	// line 1718, 1920
	wire CARRY17181920_0, CARRY17181920_1, CARRY17181920_2, CARRY17181920_3, CARRY17181920_4;
	cla l2_40(.A(W1718[3:0]), .B(W1920[3:0]), .CIN(1'b0), .COUT(CARRY17181920_0), .S(OUT17181920[3:0]));
	cla l2_41(.A(W1718[7:4]), .B(W1920[7:4]), .CIN(CARRY17181920_0), .COUT(CARRY17181920_1), .S(OUT17181920[7:4]));
	cla l2_42(.A(W1718[11:8]), .B(W1920[11:8]), .CIN(CARRY17181920_1), .COUT(CARRY17181920_2), .S(OUT17181920[11:8]));
	cla l2_43(.A(W1718[15:12]), .B(W1920[15:12]), .CIN(CARRY17181920_2), .COUT(CARRY17181920_3), .S(OUT17181920[15:12]));
	cla l2_44(.A({1'b0,W1718[18:16]}), .B(W1920[19:16]), .CIN(CARRY17181920_3), .COUT(CARRY17181920_4), .S(OUT17181920[19:16]));
	ha  l2_45(.A(W1920[20]), .B(CARRY17181920_4), .COUT(OUT17181920[21]), .SUM(OUT17181920[20]));
	
	// line 2122, 2324
	wire CARRY21222324_0, CARRY21222324_1, CARRY21222324_2, CARRY21222324_3, CARRY21222324_4, CARRY21222324_5;
	cla l2_50(.A(W2122[3:0]), .B(W2324[3:0]), .CIN(1'b0), .COUT(CARRY21222324_0), .S(OUT21222324[3:0]));
	cla l2_51(.A(W2122[7:4]), .B(W2324[7:4]), .CIN(CARRY21222324_0), .COUT(CARRY21222324_1), .S(OUT21222324[7:4]));
	cla l2_52(.A(W2122[11:8]), .B(W2324[11:8]), .CIN(CARRY21222324_1), .COUT(CARRY21222324_2), .S(OUT21222324[11:8]));
	cla l2_53(.A(W2122[15:12]), .B(W2324[15:12]), .CIN(CARRY21222324_2), .COUT(CARRY21222324_3), .S(OUT21222324[15:12]));
	cla l2_54(.A(W2122[19:16]), .B(W2324[19:16]), .CIN(CARRY21222324_3), .COUT(CARRY21222324_4), .S(OUT21222324[19:16]));
	cla l2_55(.A({1'b0,W2122[22:20]}), .B(W2324[23:20]), .CIN(CARRY21222324_4), .COUT(CARRY21222324_5), .S(OUT21222324[23:20]));
	ha  l2_56(.A(W2324[24]), .B(CARRY21222324_5), .COUT(), .SUM(OUT21222324[24]));

endmodule 

