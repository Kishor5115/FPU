



module mul_l5(W12345678910111213141516,W1718192021222324,OUT);
		input  [19:0] W12345678910111213141516;
		input  [24:0] W1718192021222324;
		output [24:0] OUT;
	// line 17181920, 21222324
	wire CARRY_0, CARRY_1, CARRY_2, CARRY_3, CARRY_4, CARRY_5;
	cla  l5_00(.A(W12345678910111213141516[3:0]), .B(W1718192021222324[3:0]), .CIN(1'b0), .COUT(CARRY_0), .S(OUT[3:0]));
	cla  l5_01(.A(W12345678910111213141516[7:4]), .B(W1718192021222324[7:4]), .CIN(CARRY_0), .COUT(CARRY_1), .S(OUT[7:4]));
	cla  l5_02(.A(W12345678910111213141516[11:8]), .B(W1718192021222324[11:8]), .CIN(CARRY_1), .COUT(CARRY_2), .S(OUT[11:8]));
	cla  l5_03(.A(W12345678910111213141516[15:12]), .B(W1718192021222324[15:12]), .CIN(CARRY_2), .COUT(CARRY_3), .S(OUT[15:12]));
	cla  l5_04(.A(W12345678910111213141516[19:16]), .B(W1718192021222324[19:16]), .CIN(CARRY_3), .COUT(CARRY_4), .S(OUT[19:16]));
	ocla l5_05(.A(W1718192021222324[23:20]), .CIN(CARRY_4), .COUT(CARRY_5), .S(OUT[23:20]));
	ha   l5_06(.A(W1718192021222324[24]), .B(CARRY_5), .COUT(), .SUM(OUT[24]));
endmodule 

